-- yet to be implemented